`ifndef TYPEDEFS_H
`define TYPEDEFS_H

package TYPEDEFS_P;

typedef logic	bool;
typedef logic[7:0] 		uint8_t;
typedef logic[15:0] 	uint16_t;
typedef logic[31:0] 	uint32_t;
typedef logic[63:0] 	uint64_t;

endpackage

`endif